module adderfp();

endmodule
